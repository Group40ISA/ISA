library verilog;
use verilog.vl_types.all;
entity tb_fp is
end tb_fp;
