library verilog;
use verilog.vl_types.all;
entity tb_uP is
end tb_uP;
